// Renan Chaves Bezerra - 121110071
// Roteiro 1

parameter divide_by=100000000;  // divisor do clock de referência
// A frequencia do clock de referencia é 50 MHz.
// A frequencia de clk_2 será de  50 MHz / divide_by

parameter NBITS_INSTR = 32;
parameter NBITS_TOP = 8, NREGS_TOP = 32, NBITS_LCD = 64;
module top(input  logic clk_2,
           input  logic [NBITS_TOP-1:0] SWI,
           output logic [NBITS_TOP-1:0] LED,
           output logic [NBITS_TOP-1:0] SEG,
           output logic [NBITS_LCD-1:0] lcd_a, lcd_b,
           output logic [NBITS_INSTR-1:0] lcd_instruction,
           output logic [NBITS_TOP-1:0] lcd_registrador [0:NREGS_TOP-1],
           output logic [NBITS_TOP-1:0] lcd_pc, lcd_SrcA, lcd_SrcB,
             lcd_ALUResult, lcd_Result, lcd_WriteData, lcd_ReadData, 
           output logic lcd_MemWrite, lcd_Branch, lcd_MemtoReg, lcd_RegWrite);

  always_comb begin
    //SEG <= SWI;
    lcd_WriteData <= SWI;
    lcd_pc <= 'h12;
    lcd_instruction <= 'h34567890;
    lcd_SrcA <= 'hab;
    lcd_SrcB <= 'hcd;
    lcd_ALUResult <= 'hef;
    lcd_Result <= 'h11;
    lcd_ReadData <= 'h33;
    lcd_MemWrite <= SWI[0];
    lcd_Branch <= SWI[1];
    lcd_MemtoReg <= SWI[2];
    lcd_RegWrite <= SWI[3];
    for(int i=0; i<NREGS_TOP; i++)
       if(i != NREGS_TOP/2-1) lcd_registrador[i] <= i+i*16;
       else                   lcd_registrador[i] <= ~SWI;
    lcd_a <= {56'h1234567890ABCD, SWI};
    lcd_b <= {SWI, 56'hFEDCBA09876543};
  end

	// COFRE
	
	logic cofre;
	logic relogio;
	logic gerente;
	logic alarme;
	
  always_comb begin
  	cofre <= SWI[0];
  	relogio <= SWI[1];
  	gerente <= SWI[2];
  end
  
  
  always_comb 
  	alarme <= cofre & (~relogio | gerente);
  
  always_comb
  	LED[1] <= alarme;
 	
  // ESTUFA
  
  logic t1;
  logic t2;
  logic a;
  logic r;
  logic i;
  
  always_comb begin
  	t1 <= SWI[7];
  	t2 <= SWI[6];
	end
	
	always_comb begin
		if (t1)
			if (t2) begin
				a <= 0;
				r <= 1;
				i <= 0;
			end
				
			else begin
				a <= 0;
				r <= 0;
				i <= 0;
				end
				
		else
			if (t2) begin
				a <= 0;
				r <= 0;
				i <= 1;
				end
				
			else begin
				a <= 1;
				r <= 0;
				i <= 0;
				end
	end
	
	always_comb begin
		LED[7] <= a;
		LED[6] <= r;
		SEG[7] <= i;
	end
	
endmodule
